//cos function lookup table
//full precision and [0 .. 45) degrees
`timescale 1ns/10ps

module cos(
    input cos_en,
    input [11:0] angle, //full angle
    output reg [15:0] result
);

reg except;
reg [14:0] cos_mem [512:0];
reg [14:0] sin_mem [512:0];
reg [9:0] angle_mem; //memory address

//logic variables
reg select_cos_mem;
reg select_positive;
reg [11:0] angle_output, angle_mem_full;
reg [14:0] mem_val;

initial begin
    //defaults
    result = 16'b0000_0000_0000_0000;
    mem_val = 15'b000_0000_0000_0000;
    angle_output = 12'b0000_0000_0000;
    angle_mem_full = 12'b0000_0000_0000;
    select_cos_mem = 1'b0;
    select_positive = 1'b1;
    //load values to memory
    cos_mem[10'b0000000000] = 15'b000000000000000; sin_mem[10'b0000000000] = 15'b000000000000000
    cos_mem[10'b0000000001] = 15'b000000000000000; sin_mem[10'b0000000001] = 15'b000000000011001
    cos_mem[10'b0000000010] = 15'b000000000000000; sin_mem[10'b0000000010] = 15'b000000000110010
    cos_mem[10'b0000000011] = 15'b000000000000000; sin_mem[10'b0000000011] = 15'b000000001001011
    cos_mem[10'b0000000100] = 15'b000000000000000; sin_mem[10'b0000000100] = 15'b000000001100101
    cos_mem[10'b0000000101] = 15'b000000000000000; sin_mem[10'b0000000101] = 15'b000000001111110
    cos_mem[10'b0000000110] = 15'b011111111111111; sin_mem[10'b0000000110] = 15'b000000010010111
    cos_mem[10'b0000000111] = 15'b011111111111111; sin_mem[10'b0000000111] = 15'b000000010110000
    cos_mem[10'b0000001000] = 15'b011111111111111; sin_mem[10'b0000001000] = 15'b000000011001001
    cos_mem[10'b0000001001] = 15'b011111111111110; sin_mem[10'b0000001001] = 15'b000000011100010
    cos_mem[10'b0000001010] = 15'b011111111111110; sin_mem[10'b0000001010] = 15'b000000011111011
    cos_mem[10'b0000001011] = 15'b011111111111110; sin_mem[10'b0000001011] = 15'b000000100010100
    cos_mem[10'b0000001100] = 15'b011111111111101; sin_mem[10'b0000001100] = 15'b000000100101110
    cos_mem[10'b0000001101] = 15'b011111111111101; sin_mem[10'b0000001101] = 15'b000000101000111
    cos_mem[10'b0000001110] = 15'b011111111111100; sin_mem[10'b0000001110] = 15'b000000101100000
//cut here -----------------------------------------------------------------------------------------
    cos_mem[10'b0000001111] = 15'b011111111111100; sin_mem[10'b0000001111] = 15'b000000101111001
    cos_mem[10'b0000010000] = 15'b011111111111011; sin_mem[10'b0000010000] = 15'b000000110010010
    cos_mem[10'b0000010001] = 15'b011111111111010; sin_mem[10'b0000010001] = 15'b000000110101011
    cos_mem[10'b0000010010] = 15'b011111111111010; sin_mem[10'b0000010010] = 15'b000000111000100
    cos_mem[10'b0000010011] = 15'b011111111111001; sin_mem[10'b0000010011] = 15'b000000111011101
    cos_mem[10'b0000010100] = 15'b011111111111000; sin_mem[10'b0000010100] = 15'b000000111110111
    cos_mem[10'b0000010101] = 15'b011111111110111; sin_mem[10'b0000010101] = 15'b000001000010000
    cos_mem[10'b0000010110] = 15'b011111111110111; sin_mem[10'b0000010110] = 15'b000001000101001
    cos_mem[10'b0000010111] = 15'b011111111110110; sin_mem[10'b0000010111] = 15'b000001001000010
    cos_mem[10'b0000011000] = 15'b011111111110101; sin_mem[10'b0000011000] = 15'b000001001011011
    cos_mem[10'b0000011001] = 15'b011111111110100; sin_mem[10'b0000011001] = 15'b000001001110100
    cos_mem[10'b0000011010] = 15'b011111111110011; sin_mem[10'b0000011010] = 15'b000001010001101
    cos_mem[10'b0000011011] = 15'b011111111110010; sin_mem[10'b0000011011] = 15'b000001010100110
    cos_mem[10'b0000011100] = 15'b011111111110001; sin_mem[10'b0000011100] = 15'b000001011000000
    cos_mem[10'b0000011101] = 15'b011111111110000; sin_mem[10'b0000011101] = 15'b000001011011001
    cos_mem[10'b0000011110] = 15'b011111111101111; sin_mem[10'b0000011110] = 15'b000001011110010
    cos_mem[10'b0000011111] = 15'b011111111101101; sin_mem[10'b0000011111] = 15'b000001100001011
    cos_mem[10'b0000100000] = 15'b011111111101100; sin_mem[10'b0000100000] = 15'b000001100100100
    cos_mem[10'b0000100001] = 15'b011111111101011; sin_mem[10'b0000100001] = 15'b000001100111101
    cos_mem[10'b0000100010] = 15'b011111111101010; sin_mem[10'b0000100010] = 15'b000001101010110
    cos_mem[10'b0000100011] = 15'b011111111101000; sin_mem[10'b0000100011] = 15'b000001101101111
    cos_mem[10'b0000100100] = 15'b011111111100111; sin_mem[10'b0000100100] = 15'b000001110001000
    cos_mem[10'b0000100101] = 15'b011111111100110; sin_mem[10'b0000100101] = 15'b000001110100001
    cos_mem[10'b0000100110] = 15'b011111111100100; sin_mem[10'b0000100110] = 15'b000001110111011
    cos_mem[10'b0000100111] = 15'b011111111100011; sin_mem[10'b0000100111] = 15'b000001111010100
    cos_mem[10'b0000101000] = 15'b011111111100001; sin_mem[10'b0000101000] = 15'b000001111101101
    cos_mem[10'b0000101001] = 15'b011111111100000; sin_mem[10'b0000101001] = 15'b000010000000110
    cos_mem[10'b0000101010] = 15'b011111111011110; sin_mem[10'b0000101010] = 15'b000010000011111
    cos_mem[10'b0000101011] = 15'b011111111011100; sin_mem[10'b0000101011] = 15'b000010000111000
    cos_mem[10'b0000101100] = 15'b011111111011011; sin_mem[10'b0000101100] = 15'b000010001010001
    cos_mem[10'b0000101101] = 15'b011111111011001; sin_mem[10'b0000101101] = 15'b000010001101010
    cos_mem[10'b0000101110] = 15'b011111111010111; sin_mem[10'b0000101110] = 15'b000010010000011
    cos_mem[10'b0000101111] = 15'b011111111010101; sin_mem[10'b0000101111] = 15'b000010010011100
    cos_mem[10'b0000110000] = 15'b011111111010100; sin_mem[10'b0000110000] = 15'b000010010110101
    cos_mem[10'b0000110001] = 15'b011111111010010; sin_mem[10'b0000110001] = 15'b000010011001110
    cos_mem[10'b0000110010] = 15'b011111111010000; sin_mem[10'b0000110010] = 15'b000010011100111
    cos_mem[10'b0000110011] = 15'b011111111001110; sin_mem[10'b0000110011] = 15'b000010100000000
    cos_mem[10'b0000110100] = 15'b011111111001100; sin_mem[10'b0000110100] = 15'b000010100011010
    cos_mem[10'b0000110101] = 15'b011111111001010; sin_mem[10'b0000110101] = 15'b000010100110011
    cos_mem[10'b0000110110] = 15'b011111111001000; sin_mem[10'b0000110110] = 15'b000010101001100
    cos_mem[10'b0000110111] = 15'b011111111000110; sin_mem[10'b0000110111] = 15'b000010101100101
    cos_mem[10'b0000111000] = 15'b011111111000100; sin_mem[10'b0000111000] = 15'b000010101111110
    cos_mem[10'b0000111001] = 15'b011111111000001; sin_mem[10'b0000111001] = 15'b000010110010111
    cos_mem[10'b0000111010] = 15'b011111110111111; sin_mem[10'b0000111010] = 15'b000010110110000
    cos_mem[10'b0000111011] = 15'b011111110111101; sin_mem[10'b0000111011] = 15'b000010111001001
    cos_mem[10'b0000111100] = 15'b011111110111011; sin_mem[10'b0000111100] = 15'b000010111100010
    cos_mem[10'b0000111101] = 15'b011111110111000; sin_mem[10'b0000111101] = 15'b000010111111011
    cos_mem[10'b0000111110] = 15'b011111110110110; sin_mem[10'b0000111110] = 15'b000011000010100
    cos_mem[10'b0000111111] = 15'b011111110110100; sin_mem[10'b0000111111] = 15'b000011000101101
    cos_mem[10'b0001000000] = 15'b011111110110001; sin_mem[10'b0001000000] = 15'b000011001000110
    cos_mem[10'b0001000001] = 15'b011111110101111; sin_mem[10'b0001000001] = 15'b000011001011111
    cos_mem[10'b0001000010] = 15'b011111110101100; sin_mem[10'b0001000010] = 15'b000011001111000
    cos_mem[10'b0001000011] = 15'b011111110101010; sin_mem[10'b0001000011] = 15'b000011010010001
    cos_mem[10'b0001000100] = 15'b011111110100111; sin_mem[10'b0001000100] = 15'b000011010101010
    cos_mem[10'b0001000101] = 15'b011111110100100; sin_mem[10'b0001000101] = 15'b000011011000011
    cos_mem[10'b0001000110] = 15'b011111110100010; sin_mem[10'b0001000110] = 15'b000011011011100
    cos_mem[10'b0001000111] = 15'b011111110011111; sin_mem[10'b0001000111] = 15'b000011011110101
    cos_mem[10'b0001001000] = 15'b011111110011100; sin_mem[10'b0001001000] = 15'b000011100001110
    cos_mem[10'b0001001001] = 15'b011111110011001; sin_mem[10'b0001001001] = 15'b000011100100111
    cos_mem[10'b0001001010] = 15'b011111110010111; sin_mem[10'b0001001010] = 15'b000011101000000
    cos_mem[10'b0001001011] = 15'b011111110010100; sin_mem[10'b0001001011] = 15'b000011101011001
    cos_mem[10'b0001001100] = 15'b011111110010001; sin_mem[10'b0001001100] = 15'b000011101110010
    cos_mem[10'b0001001101] = 15'b011111110001110; sin_mem[10'b0001001101] = 15'b000011110001011
    cos_mem[10'b0001001110] = 15'b011111110001011; sin_mem[10'b0001001110] = 15'b000011110100100
    cos_mem[10'b0001001111] = 15'b011111110001000; sin_mem[10'b0001001111] = 15'b000011110111101
    cos_mem[10'b0001010000] = 15'b011111110000101; sin_mem[10'b0001010000] = 15'b000011111010110
    cos_mem[10'b0001010001] = 15'b011111110000010; sin_mem[10'b0001010001] = 15'b000011111101111
    cos_mem[10'b0001010010] = 15'b011111101111111; sin_mem[10'b0001010010] = 15'b000100000000111
    cos_mem[10'b0001010011] = 15'b011111101111011; sin_mem[10'b0001010011] = 15'b000100000100000
    cos_mem[10'b0001010100] = 15'b011111101111000; sin_mem[10'b0001010100] = 15'b000100000111001
    cos_mem[10'b0001010101] = 15'b011111101110101; sin_mem[10'b0001010101] = 15'b000100001010010
    cos_mem[10'b0001010110] = 15'b011111101110010; sin_mem[10'b0001010110] = 15'b000100001101011
    cos_mem[10'b0001010111] = 15'b011111101101110; sin_mem[10'b0001010111] = 15'b000100010000100
    cos_mem[10'b0001011000] = 15'b011111101101011; sin_mem[10'b0001011000] = 15'b000100010011101
    cos_mem[10'b0001011001] = 15'b011111101101000; sin_mem[10'b0001011001] = 15'b000100010110110
    cos_mem[10'b0001011010] = 15'b011111101100100; sin_mem[10'b0001011010] = 15'b000100011001111
    cos_mem[10'b0001011011] = 15'b011111101100001; sin_mem[10'b0001011011] = 15'b000100011101000
    cos_mem[10'b0001011100] = 15'b011111101011101; sin_mem[10'b0001011100] = 15'b000100100000001
    cos_mem[10'b0001011101] = 15'b011111101011010; sin_mem[10'b0001011101] = 15'b000100100011001
    cos_mem[10'b0001011110] = 15'b011111101010110; sin_mem[10'b0001011110] = 15'b000100100110010
    cos_mem[10'b0001011111] = 15'b011111101010010; sin_mem[10'b0001011111] = 15'b000100101001011
    cos_mem[10'b0001100000] = 15'b011111101001111; sin_mem[10'b0001100000] = 15'b000100101100100
    cos_mem[10'b0001100001] = 15'b011111101001011; sin_mem[10'b0001100001] = 15'b000100101111101
    cos_mem[10'b0001100010] = 15'b011111101000111; sin_mem[10'b0001100010] = 15'b000100110010110
    cos_mem[10'b0001100011] = 15'b011111101000011; sin_mem[10'b0001100011] = 15'b000100110101111
    cos_mem[10'b0001100100] = 15'b011111101000000; sin_mem[10'b0001100100] = 15'b000100111000111
    cos_mem[10'b0001100101] = 15'b011111100111100; sin_mem[10'b0001100101] = 15'b000100111100000
    cos_mem[10'b0001100110] = 15'b011111100111000; sin_mem[10'b0001100110] = 15'b000100111111001
    cos_mem[10'b0001100111] = 15'b011111100110100; sin_mem[10'b0001100111] = 15'b000101000010010
    cos_mem[10'b0001101000] = 15'b011111100110000; sin_mem[10'b0001101000] = 15'b000101000101011
    cos_mem[10'b0001101001] = 15'b011111100101100; sin_mem[10'b0001101001] = 15'b000101001000100
    cos_mem[10'b0001101010] = 15'b011111100101000; sin_mem[10'b0001101010] = 15'b000101001011100
    cos_mem[10'b0001101011] = 15'b011111100100100; sin_mem[10'b0001101011] = 15'b000101001110101
    cos_mem[10'b0001101100] = 15'b011111100100000; sin_mem[10'b0001101100] = 15'b000101010001110
    cos_mem[10'b0001101101] = 15'b011111100011100; sin_mem[10'b0001101101] = 15'b000101010100111
    cos_mem[10'b0001101110] = 15'b011111100010111; sin_mem[10'b0001101110] = 15'b000101011000000
    cos_mem[10'b0001101111] = 15'b011111100010011; sin_mem[10'b0001101111] = 15'b000101011011000
    cos_mem[10'b0001110000] = 15'b011111100001111; sin_mem[10'b0001110000] = 15'b000101011110001
    cos_mem[10'b0001110001] = 15'b011111100001010; sin_mem[10'b0001110001] = 15'b000101100001010
    cos_mem[10'b0001110010] = 15'b011111100000110; sin_mem[10'b0001110010] = 15'b000101100100011
    cos_mem[10'b0001110011] = 15'b011111100000010; sin_mem[10'b0001110011] = 15'b000101100111011
    cos_mem[10'b0001110100] = 15'b011111011111101; sin_mem[10'b0001110100] = 15'b000101101010100
    cos_mem[10'b0001110101] = 15'b011111011111001; sin_mem[10'b0001110101] = 15'b000101101101101
    cos_mem[10'b0001110110] = 15'b011111011110100; sin_mem[10'b0001110110] = 15'b000101110000101
    cos_mem[10'b0001110111] = 15'b011111011110000; sin_mem[10'b0001110111] = 15'b000101110011110
    cos_mem[10'b0001111000] = 15'b011111011101011; sin_mem[10'b0001111000] = 15'b000101110110111
    cos_mem[10'b0001111001] = 15'b011111011100111; sin_mem[10'b0001111001] = 15'b000101111010000
    cos_mem[10'b0001111010] = 15'b011111011100010; sin_mem[10'b0001111010] = 15'b000101111101000
    cos_mem[10'b0001111011] = 15'b011111011011101; sin_mem[10'b0001111011] = 15'b000110000000001
    cos_mem[10'b0001111100] = 15'b011111011011000; sin_mem[10'b0001111100] = 15'b000110000011010
    cos_mem[10'b0001111101] = 15'b011111011010100; sin_mem[10'b0001111101] = 15'b000110000110010
    cos_mem[10'b0001111110] = 15'b011111011001111; sin_mem[10'b0001111110] = 15'b000110001001011
    cos_mem[10'b0001111111] = 15'b011111011001010; sin_mem[10'b0001111111] = 15'b000110001100100
    cos_mem[10'b0010000000] = 15'b011111011000101; sin_mem[10'b0010000000] = 15'b000110001111100
    cos_mem[10'b0010000001] = 15'b011111011000000; sin_mem[10'b0010000001] = 15'b000110010010101
    cos_mem[10'b0010000010] = 15'b011111010111011; sin_mem[10'b0010000010] = 15'b000110010101110
    cos_mem[10'b0010000011] = 15'b011111010110110; sin_mem[10'b0010000011] = 15'b000110011000110
    cos_mem[10'b0010000100] = 15'b011111010110001; sin_mem[10'b0010000100] = 15'b000110011011111
    cos_mem[10'b0010000101] = 15'b011111010101100; sin_mem[10'b0010000101] = 15'b000110011111000
    cos_mem[10'b0010000110] = 15'b011111010100111; sin_mem[10'b0010000110] = 15'b000110100010000
    cos_mem[10'b0010000111] = 15'b011111010100010; sin_mem[10'b0010000111] = 15'b000110100101001
    cos_mem[10'b0010001000] = 15'b011111010011101; sin_mem[10'b0010001000] = 15'b000110101000001
    cos_mem[10'b0010001001] = 15'b011111010011000; sin_mem[10'b0010001001] = 15'b000110101011010
    cos_mem[10'b0010001010] = 15'b011111010010010; sin_mem[10'b0010001010] = 15'b000110101110010
    cos_mem[10'b0010001011] = 15'b011111010001101; sin_mem[10'b0010001011] = 15'b000110110001011
    cos_mem[10'b0010001100] = 15'b011111010001000; sin_mem[10'b0010001100] = 15'b000110110100100
    cos_mem[10'b0010001101] = 15'b011111010000010; sin_mem[10'b0010001101] = 15'b000110110111100
    cos_mem[10'b0010001110] = 15'b011111001111101; sin_mem[10'b0010001110] = 15'b000110111010101
    cos_mem[10'b0010001111] = 15'b011111001110111; sin_mem[10'b0010001111] = 15'b000110111101101
    cos_mem[10'b0010010000] = 15'b011111001110010; sin_mem[10'b0010010000] = 15'b000111000000110
    cos_mem[10'b0010010001] = 15'b011111001101100; sin_mem[10'b0010010001] = 15'b000111000011110
    cos_mem[10'b0010010010] = 15'b011111001100111; sin_mem[10'b0010010010] = 15'b000111000110111
    cos_mem[10'b0010010011] = 15'b011111001100001; sin_mem[10'b0010010011] = 15'b000111001001111
    cos_mem[10'b0010010100] = 15'b011111001011100; sin_mem[10'b0010010100] = 15'b000111001101000
    cos_mem[10'b0010010101] = 15'b011111001010110; sin_mem[10'b0010010101] = 15'b000111010000000
    cos_mem[10'b0010010110] = 15'b011111001010000; sin_mem[10'b0010010110] = 15'b000111010011001
    cos_mem[10'b0010010111] = 15'b011111001001010; sin_mem[10'b0010010111] = 15'b000111010110001
    cos_mem[10'b0010011000] = 15'b011111001000101; sin_mem[10'b0010011000] = 15'b000111011001010
    cos_mem[10'b0010011001] = 15'b011111000111111; sin_mem[10'b0010011001] = 15'b000111011100010
    cos_mem[10'b0010011010] = 15'b011111000111001; sin_mem[10'b0010011010] = 15'b000111011111011
    cos_mem[10'b0010011011] = 15'b011111000110011; sin_mem[10'b0010011011] = 15'b000111100010011
    cos_mem[10'b0010011100] = 15'b011111000101101; sin_mem[10'b0010011100] = 15'b000111100101011
    cos_mem[10'b0010011101] = 15'b011111000100111; sin_mem[10'b0010011101] = 15'b000111101000100
    cos_mem[10'b0010011110] = 15'b011111000100001; sin_mem[10'b0010011110] = 15'b000111101011100
    cos_mem[10'b0010011111] = 15'b011111000011011; sin_mem[10'b0010011111] = 15'b000111101110101
    cos_mem[10'b0010100000] = 15'b011111000010101; sin_mem[10'b0010100000] = 15'b000111110001101
    cos_mem[10'b0010100001] = 15'b011111000001111; sin_mem[10'b0010100001] = 15'b000111110100101
    cos_mem[10'b0010100010] = 15'b011111000001001; sin_mem[10'b0010100010] = 15'b000111110111110
    cos_mem[10'b0010100011] = 15'b011111000000011; sin_mem[10'b0010100011] = 15'b000111111010110
    cos_mem[10'b0010100100] = 15'b011110111111100; sin_mem[10'b0010100100] = 15'b000111111101110
    cos_mem[10'b0010100101] = 15'b011110111110110; sin_mem[10'b0010100101] = 15'b001000000000111
    cos_mem[10'b0010100110] = 15'b011110111110000; sin_mem[10'b0010100110] = 15'b001000000011111
    cos_mem[10'b0010100111] = 15'b011110111101001; sin_mem[10'b0010100111] = 15'b001000000110111
    cos_mem[10'b0010101000] = 15'b011110111100011; sin_mem[10'b0010101000] = 15'b001000001010000
    cos_mem[10'b0010101001] = 15'b011110111011101; sin_mem[10'b0010101001] = 15'b001000001101000
    cos_mem[10'b0010101010] = 15'b011110111010110; sin_mem[10'b0010101010] = 15'b001000010000000
    cos_mem[10'b0010101011] = 15'b011110111010000; sin_mem[10'b0010101011] = 15'b001000010011001
    cos_mem[10'b0010101100] = 15'b011110111001001; sin_mem[10'b0010101100] = 15'b001000010110001
    cos_mem[10'b0010101101] = 15'b011110111000010; sin_mem[10'b0010101101] = 15'b001000011001001
    cos_mem[10'b0010101110] = 15'b011110110111100; sin_mem[10'b0010101110] = 15'b001000011100001
    cos_mem[10'b0010101111] = 15'b011110110110101; sin_mem[10'b0010101111] = 15'b001000011111010
    cos_mem[10'b0010110000] = 15'b011110110101111; sin_mem[10'b0010110000] = 15'b001000100010010
    cos_mem[10'b0010110001] = 15'b011110110101000; sin_mem[10'b0010110001] = 15'b001000100101010
    cos_mem[10'b0010110010] = 15'b011110110100001; sin_mem[10'b0010110010] = 15'b001000101000010
    cos_mem[10'b0010110011] = 15'b011110110011010; sin_mem[10'b0010110011] = 15'b001000101011010
    cos_mem[10'b0010110100] = 15'b011110110010011; sin_mem[10'b0010110100] = 15'b001000101110011
    cos_mem[10'b0010110101] = 15'b011110110001101; sin_mem[10'b0010110101] = 15'b001000110001011
    cos_mem[10'b0010110110] = 15'b011110110000110; sin_mem[10'b0010110110] = 15'b001000110100011
    cos_mem[10'b0010110111] = 15'b011110101111111; sin_mem[10'b0010110111] = 15'b001000110111011
    cos_mem[10'b0010111000] = 15'b011110101111000; sin_mem[10'b0010111000] = 15'b001000111010011
    cos_mem[10'b0010111001] = 15'b011110101110001; sin_mem[10'b0010111001] = 15'b001000111101011
    cos_mem[10'b0010111010] = 15'b011110101101010; sin_mem[10'b0010111010] = 15'b001001000000100
    cos_mem[10'b0010111011] = 15'b011110101100011; sin_mem[10'b0010111011] = 15'b001001000011100
    cos_mem[10'b0010111100] = 15'b011110101011011; sin_mem[10'b0010111100] = 15'b001001000110100
    cos_mem[10'b0010111101] = 15'b011110101010100; sin_mem[10'b0010111101] = 15'b001001001001100
    cos_mem[10'b0010111110] = 15'b011110101001101; sin_mem[10'b0010111110] = 15'b001001001100100
    cos_mem[10'b0010111111] = 15'b011110101000110; sin_mem[10'b0010111111] = 15'b001001001111100
    cos_mem[10'b0011000000] = 15'b011110100111111; sin_mem[10'b0011000000] = 15'b001001010010100
    cos_mem[10'b0011000001] = 15'b011110100110111; sin_mem[10'b0011000001] = 15'b001001010101100
    cos_mem[10'b0011000010] = 15'b011110100110000; sin_mem[10'b0011000010] = 15'b001001011000100
    cos_mem[10'b0011000011] = 15'b011110100101000; sin_mem[10'b0011000011] = 15'b001001011011100
    cos_mem[10'b0011000100] = 15'b011110100100001; sin_mem[10'b0011000100] = 15'b001001011110100
    cos_mem[10'b0011000101] = 15'b011110100011010; sin_mem[10'b0011000101] = 15'b001001100001100
    cos_mem[10'b0011000110] = 15'b011110100010010; sin_mem[10'b0011000110] = 15'b001001100100100
    cos_mem[10'b0011000111] = 15'b011110100001011; sin_mem[10'b0011000111] = 15'b001001100111100
    cos_mem[10'b0011001000] = 15'b011110100000011; sin_mem[10'b0011001000] = 15'b001001101010100
    cos_mem[10'b0011001001] = 15'b011110011111011; sin_mem[10'b0011001001] = 15'b001001101101100
    cos_mem[10'b0011001010] = 15'b011110011110100; sin_mem[10'b0011001010] = 15'b001001110000100
    cos_mem[10'b0011001011] = 15'b011110011101100; sin_mem[10'b0011001011] = 15'b001001110011100
    cos_mem[10'b0011001100] = 15'b011110011100100; sin_mem[10'b0011001100] = 15'b001001110110100
    cos_mem[10'b0011001101] = 15'b011110011011101; sin_mem[10'b0011001101] = 15'b001001111001100
    cos_mem[10'b0011001110] = 15'b011110011010101; sin_mem[10'b0011001110] = 15'b001001111100100
    cos_mem[10'b0011001111] = 15'b011110011001101; sin_mem[10'b0011001111] = 15'b001001111111011
    cos_mem[10'b0011010000] = 15'b011110011000101; sin_mem[10'b0011010000] = 15'b001010000010011
    cos_mem[10'b0011010001] = 15'b011110010111101; sin_mem[10'b0011010001] = 15'b001010000101011
    cos_mem[10'b0011010010] = 15'b011110010110101; sin_mem[10'b0011010010] = 15'b001010001000011
    cos_mem[10'b0011010011] = 15'b011110010101101; sin_mem[10'b0011010011] = 15'b001010001011011
    cos_mem[10'b0011010100] = 15'b011110010100101; sin_mem[10'b0011010100] = 15'b001010001110011
    cos_mem[10'b0011010101] = 15'b011110010011101; sin_mem[10'b0011010101] = 15'b001010010001011
    cos_mem[10'b0011010110] = 15'b011110010010101; sin_mem[10'b0011010110] = 15'b001010010100010
    cos_mem[10'b0011010111] = 15'b011110010001101; sin_mem[10'b0011010111] = 15'b001010010111010
    cos_mem[10'b0011011000] = 15'b011110010000101; sin_mem[10'b0011011000] = 15'b001010011010010
    cos_mem[10'b0011011001] = 15'b011110001111101; sin_mem[10'b0011011001] = 15'b001010011101010
    cos_mem[10'b0011011010] = 15'b011110001110100; sin_mem[10'b0011011010] = 15'b001010100000001
    cos_mem[10'b0011011011] = 15'b011110001101100; sin_mem[10'b0011011011] = 15'b001010100011001
    cos_mem[10'b0011011100] = 15'b011110001100100; sin_mem[10'b0011011100] = 15'b001010100110001
    cos_mem[10'b0011011101] = 15'b011110001011011; sin_mem[10'b0011011101] = 15'b001010101001001
    cos_mem[10'b0011011110] = 15'b011110001010011; sin_mem[10'b0011011110] = 15'b001010101100000
    cos_mem[10'b0011011111] = 15'b011110001001011; sin_mem[10'b0011011111] = 15'b001010101111000
    cos_mem[10'b0011100000] = 15'b011110001000010; sin_mem[10'b0011100000] = 15'b001010110010000
    cos_mem[10'b0011100001] = 15'b011110000111010; sin_mem[10'b0011100001] = 15'b001010110100111
    cos_mem[10'b0011100010] = 15'b011110000110001; sin_mem[10'b0011100010] = 15'b001010110111111
    cos_mem[10'b0011100011] = 15'b011110000101001; sin_mem[10'b0011100011] = 15'b001010111010111
    cos_mem[10'b0011100100] = 15'b011110000100000; sin_mem[10'b0011100100] = 15'b001010111101110
    cos_mem[10'b0011100101] = 15'b011110000010111; sin_mem[10'b0011100101] = 15'b001011000000110
    cos_mem[10'b0011100110] = 15'b011110000001111; sin_mem[10'b0011100110] = 15'b001011000011101
    cos_mem[10'b0011100111] = 15'b011110000000110; sin_mem[10'b0011100111] = 15'b001011000110101
    cos_mem[10'b0011101000] = 15'b011101111111101; sin_mem[10'b0011101000] = 15'b001011001001100
    cos_mem[10'b0011101001] = 15'b011101111110101; sin_mem[10'b0011101001] = 15'b001011001100100
    cos_mem[10'b0011101010] = 15'b011101111101100; sin_mem[10'b0011101010] = 15'b001011001111100
    cos_mem[10'b0011101011] = 15'b011101111100011; sin_mem[10'b0011101011] = 15'b001011010010011
    cos_mem[10'b0011101100] = 15'b011101111011010; sin_mem[10'b0011101100] = 15'b001011010101011
    cos_mem[10'b0011101101] = 15'b011101111010001; sin_mem[10'b0011101101] = 15'b001011011000010
    cos_mem[10'b0011101110] = 15'b011101111001000; sin_mem[10'b0011101110] = 15'b001011011011010
    cos_mem[10'b0011101111] = 15'b011101110111111; sin_mem[10'b0011101111] = 15'b001011011110001
    cos_mem[10'b0011110000] = 15'b011101110110110; sin_mem[10'b0011110000] = 15'b001011100001001
    cos_mem[10'b0011110001] = 15'b011101110101101; sin_mem[10'b0011110001] = 15'b001011100100000
    cos_mem[10'b0011110010] = 15'b011101110100100; sin_mem[10'b0011110010] = 15'b001011100110111
    cos_mem[10'b0011110011] = 15'b011101110011011; sin_mem[10'b0011110011] = 15'b001011101001111
    cos_mem[10'b0011110100] = 15'b011101110010010; sin_mem[10'b0011110100] = 15'b001011101100110
    cos_mem[10'b0011110101] = 15'b011101110001000; sin_mem[10'b0011110101] = 15'b001011101111110
    cos_mem[10'b0011110110] = 15'b011101101111111; sin_mem[10'b0011110110] = 15'b001011110010101
    cos_mem[10'b0011110111] = 15'b011101101110110; sin_mem[10'b0011110111] = 15'b001011110101100
    cos_mem[10'b0011111000] = 15'b011101101101101; sin_mem[10'b0011111000] = 15'b001011111000100
    cos_mem[10'b0011111001] = 15'b011101101100011; sin_mem[10'b0011111001] = 15'b001011111011011
    cos_mem[10'b0011111010] = 15'b011101101011010; sin_mem[10'b0011111010] = 15'b001011111110010
    cos_mem[10'b0011111011] = 15'b011101101010000; sin_mem[10'b0011111011] = 15'b001100000001010
    cos_mem[10'b0011111100] = 15'b011101101000111; sin_mem[10'b0011111100] = 15'b001100000100001
    cos_mem[10'b0011111101] = 15'b011101100111110; sin_mem[10'b0011111101] = 15'b001100000111000
    cos_mem[10'b0011111110] = 15'b011101100110100; sin_mem[10'b0011111110] = 15'b001100001001111
    cos_mem[10'b0011111111] = 15'b011101100101010; sin_mem[10'b0011111111] = 15'b001100001100111
    cos_mem[10'b0100000000] = 15'b011101100100001; sin_mem[10'b0100000000] = 15'b001100001111110
    cos_mem[10'b0100000001] = 15'b011101100010111; sin_mem[10'b0100000001] = 15'b001100010010101
    cos_mem[10'b0100000010] = 15'b011101100001110; sin_mem[10'b0100000010] = 15'b001100010101100
    cos_mem[10'b0100000011] = 15'b011101100000100; sin_mem[10'b0100000011] = 15'b001100011000011
    cos_mem[10'b0100000100] = 15'b011101011111010; sin_mem[10'b0100000100] = 15'b001100011011011
    cos_mem[10'b0100000101] = 15'b011101011110000; sin_mem[10'b0100000101] = 15'b001100011110010
    cos_mem[10'b0100000110] = 15'b011101011100110; sin_mem[10'b0100000110] = 15'b001100100001001
    cos_mem[10'b0100000111] = 15'b011101011011101; sin_mem[10'b0100000111] = 15'b001100100100000
    cos_mem[10'b0100001000] = 15'b011101011010011; sin_mem[10'b0100001000] = 15'b001100100110111
    cos_mem[10'b0100001001] = 15'b011101011001001; sin_mem[10'b0100001001] = 15'b001100101001110
    cos_mem[10'b0100001010] = 15'b011101010111111; sin_mem[10'b0100001010] = 15'b001100101100101
    cos_mem[10'b0100001011] = 15'b011101010110101; sin_mem[10'b0100001011] = 15'b001100101111100
    cos_mem[10'b0100001100] = 15'b011101010101011; sin_mem[10'b0100001100] = 15'b001100110010011
    cos_mem[10'b0100001101] = 15'b011101010100001; sin_mem[10'b0100001101] = 15'b001100110101010
    cos_mem[10'b0100001110] = 15'b011101010010111; sin_mem[10'b0100001110] = 15'b001100111000001
    cos_mem[10'b0100001111] = 15'b011101010001101; sin_mem[10'b0100001111] = 15'b001100111011000
    cos_mem[10'b0100010000] = 15'b011101010000010; sin_mem[10'b0100010000] = 15'b001100111101111
    cos_mem[10'b0100010001] = 15'b011101001111000; sin_mem[10'b0100010001] = 15'b001101000000110
    cos_mem[10'b0100010010] = 15'b011101001101110; sin_mem[10'b0100010010] = 15'b001101000011101
    cos_mem[10'b0100010011] = 15'b011101001100100; sin_mem[10'b0100010011] = 15'b001101000110100
    cos_mem[10'b0100010100] = 15'b011101001011001; sin_mem[10'b0100010100] = 15'b001101001001011
    cos_mem[10'b0100010101] = 15'b011101001001111; sin_mem[10'b0100010101] = 15'b001101001100010
    cos_mem[10'b0100010110] = 15'b011101001000101; sin_mem[10'b0100010110] = 15'b001101001111001
    cos_mem[10'b0100010111] = 15'b011101000111010; sin_mem[10'b0100010111] = 15'b001101010010000
    cos_mem[10'b0100011000] = 15'b011101000110000; sin_mem[10'b0100011000] = 15'b001101010100111
    cos_mem[10'b0100011001] = 15'b011101000100101; sin_mem[10'b0100011001] = 15'b001101010111110
    cos_mem[10'b0100011010] = 15'b011101000011011; sin_mem[10'b0100011010] = 15'b001101011010100
    cos_mem[10'b0100011011] = 15'b011101000010000; sin_mem[10'b0100011011] = 15'b001101011101011
    cos_mem[10'b0100011100] = 15'b011101000000110; sin_mem[10'b0100011100] = 15'b001101100000010
    cos_mem[10'b0100011101] = 15'b011100111111011; sin_mem[10'b0100011101] = 15'b001101100011001
    cos_mem[10'b0100011110] = 15'b011100111110000; sin_mem[10'b0100011110] = 15'b001101100110000
    cos_mem[10'b0100011111] = 15'b011100111100110; sin_mem[10'b0100011111] = 15'b001101101000110
    cos_mem[10'b0100100000] = 15'b011100111011011; sin_mem[10'b0100100000] = 15'b001101101011101
    cos_mem[10'b0100100001] = 15'b011100111010000; sin_mem[10'b0100100001] = 15'b001101101110100
    cos_mem[10'b0100100010] = 15'b011100111000101; sin_mem[10'b0100100010] = 15'b001101110001010
    cos_mem[10'b0100100011] = 15'b011100110111011; sin_mem[10'b0100100011] = 15'b001101110100001
    cos_mem[10'b0100100100] = 15'b011100110110000; sin_mem[10'b0100100100] = 15'b001101110111000
    cos_mem[10'b0100100101] = 15'b011100110100101; sin_mem[10'b0100100101] = 15'b001101111001110
    cos_mem[10'b0100100110] = 15'b011100110011010; sin_mem[10'b0100100110] = 15'b001101111100101
    cos_mem[10'b0100100111] = 15'b011100110001111; sin_mem[10'b0100100111] = 15'b001101111111100
    cos_mem[10'b0100101000] = 15'b011100110000100; sin_mem[10'b0100101000] = 15'b001110000010010
    cos_mem[10'b0100101001] = 15'b011100101111001; sin_mem[10'b0100101001] = 15'b001110000101001
    cos_mem[10'b0100101010] = 15'b011100101101110; sin_mem[10'b0100101010] = 15'b001110000111111
    cos_mem[10'b0100101011] = 15'b011100101100011; sin_mem[10'b0100101011] = 15'b001110001010110
    cos_mem[10'b0100101100] = 15'b011100101011000; sin_mem[10'b0100101100] = 15'b001110001101100
    cos_mem[10'b0100101101] = 15'b011100101001100; sin_mem[10'b0100101101] = 15'b001110010000011
    cos_mem[10'b0100101110] = 15'b011100101000001; sin_mem[10'b0100101110] = 15'b001110010011001
    cos_mem[10'b0100101111] = 15'b011100100110110; sin_mem[10'b0100101111] = 15'b001110010110000
    cos_mem[10'b0100110000] = 15'b011100100101011; sin_mem[10'b0100110000] = 15'b001110011000110
    cos_mem[10'b0100110001] = 15'b011100100011111; sin_mem[10'b0100110001] = 15'b001110011011101
    cos_mem[10'b0100110010] = 15'b011100100010100; sin_mem[10'b0100110010] = 15'b001110011110011
    cos_mem[10'b0100110011] = 15'b011100100001001; sin_mem[10'b0100110011] = 15'b001110100001010
    cos_mem[10'b0100110100] = 15'b011100011111101; sin_mem[10'b0100110100] = 15'b001110100100000
    cos_mem[10'b0100110101] = 15'b011100011110010; sin_mem[10'b0100110101] = 15'b001110100110110
    cos_mem[10'b0100110110] = 15'b011100011100110; sin_mem[10'b0100110110] = 15'b001110101001101
    cos_mem[10'b0100110111] = 15'b011100011011011; sin_mem[10'b0100110111] = 15'b001110101100011
    cos_mem[10'b0100111000] = 15'b011100011001111; sin_mem[10'b0100111000] = 15'b001110101111001
    cos_mem[10'b0100111001] = 15'b011100011000011; sin_mem[10'b0100111001] = 15'b001110110010000
    cos_mem[10'b0100111010] = 15'b011100010111000; sin_mem[10'b0100111010] = 15'b001110110100110
    cos_mem[10'b0100111011] = 15'b011100010101100; sin_mem[10'b0100111011] = 15'b001110110111100
    cos_mem[10'b0100111100] = 15'b011100010100001; sin_mem[10'b0100111100] = 15'b001110111010011
    cos_mem[10'b0100111101] = 15'b011100010010101; sin_mem[10'b0100111101] = 15'b001110111101001
    cos_mem[10'b0100111110] = 15'b011100010001001; sin_mem[10'b0100111110] = 15'b001110111111111
    cos_mem[10'b0100111111] = 15'b011100001111101; sin_mem[10'b0100111111] = 15'b001111000010101
    cos_mem[10'b0101000000] = 15'b011100001110001; sin_mem[10'b0101000000] = 15'b001111000101011
    cos_mem[10'b0101000001] = 15'b011100001100110; sin_mem[10'b0101000001] = 15'b001111001000010
    cos_mem[10'b0101000010] = 15'b011100001011010; sin_mem[10'b0101000010] = 15'b001111001011000
    cos_mem[10'b0101000011] = 15'b011100001001110; sin_mem[10'b0101000011] = 15'b001111001101110
    cos_mem[10'b0101000100] = 15'b011100001000010; sin_mem[10'b0101000100] = 15'b001111010000100
    cos_mem[10'b0101000101] = 15'b011100000110110; sin_mem[10'b0101000101] = 15'b001111010011010
    cos_mem[10'b0101000110] = 15'b011100000101010; sin_mem[10'b0101000110] = 15'b001111010110000
    cos_mem[10'b0101000111] = 15'b011100000011110; sin_mem[10'b0101000111] = 15'b001111011000110
    cos_mem[10'b0101001000] = 15'b011100000010010; sin_mem[10'b0101001000] = 15'b001111011011100
    cos_mem[10'b0101001001] = 15'b011100000000101; sin_mem[10'b0101001001] = 15'b001111011110010
    cos_mem[10'b0101001010] = 15'b011011111111001; sin_mem[10'b0101001010] = 15'b001111100001000
    cos_mem[10'b0101001011] = 15'b011011111101101; sin_mem[10'b0101001011] = 15'b001111100011110
    cos_mem[10'b0101001100] = 15'b011011111100001; sin_mem[10'b0101001100] = 15'b001111100110100
    cos_mem[10'b0101001101] = 15'b011011111010101; sin_mem[10'b0101001101] = 15'b001111101001010
    cos_mem[10'b0101001110] = 15'b011011111001000; sin_mem[10'b0101001110] = 15'b001111101100000
    cos_mem[10'b0101001111] = 15'b011011110111100; sin_mem[10'b0101001111] = 15'b001111101110110
    cos_mem[10'b0101010000] = 15'b011011110110000; sin_mem[10'b0101010000] = 15'b001111110001100
    cos_mem[10'b0101010001] = 15'b011011110100011; sin_mem[10'b0101010001] = 15'b001111110100010
    cos_mem[10'b0101010010] = 15'b011011110010111; sin_mem[10'b0101010010] = 15'b001111110110111
    cos_mem[10'b0101010011] = 15'b011011110001010; sin_mem[10'b0101010011] = 15'b001111111001101
    cos_mem[10'b0101010100] = 15'b011011101111110; sin_mem[10'b0101010100] = 15'b001111111100011
    cos_mem[10'b0101010101] = 15'b011011101110001; sin_mem[10'b0101010101] = 15'b001111111111001
    cos_mem[10'b0101010110] = 15'b011011101100101; sin_mem[10'b0101010110] = 15'b010000000001111
    cos_mem[10'b0101010111] = 15'b011011101011000; sin_mem[10'b0101010111] = 15'b010000000100100
    cos_mem[10'b0101011000] = 15'b011011101001011; sin_mem[10'b0101011000] = 15'b010000000111010
    cos_mem[10'b0101011001] = 15'b011011100111111; sin_mem[10'b0101011001] = 15'b010000001010000
    cos_mem[10'b0101011010] = 15'b011011100110010; sin_mem[10'b0101011010] = 15'b010000001100101
    cos_mem[10'b0101011011] = 15'b011011100100101; sin_mem[10'b0101011011] = 15'b010000001111011
    cos_mem[10'b0101011100] = 15'b011011100011000; sin_mem[10'b0101011100] = 15'b010000010010001
    cos_mem[10'b0101011101] = 15'b011011100001100; sin_mem[10'b0101011101] = 15'b010000010100110
    cos_mem[10'b0101011110] = 15'b011011011111111; sin_mem[10'b0101011110] = 15'b010000010111100
    cos_mem[10'b0101011111] = 15'b011011011110010; sin_mem[10'b0101011111] = 15'b010000011010001
    cos_mem[10'b0101100000] = 15'b011011011100101; sin_mem[10'b0101100000] = 15'b010000011100111
    cos_mem[10'b0101100001] = 15'b011011011011000; sin_mem[10'b0101100001] = 15'b010000011111101
    cos_mem[10'b0101100010] = 15'b011011011001011; sin_mem[10'b0101100010] = 15'b010000100010010
    cos_mem[10'b0101100011] = 15'b011011010111110; sin_mem[10'b0101100011] = 15'b010000100101000
    cos_mem[10'b0101100100] = 15'b011011010110001; sin_mem[10'b0101100100] = 15'b010000100111101
    cos_mem[10'b0101100101] = 15'b011011010100100; sin_mem[10'b0101100101] = 15'b010000101010011
    cos_mem[10'b0101100110] = 15'b011011010010111; sin_mem[10'b0101100110] = 15'b010000101101000
    cos_mem[10'b0101100111] = 15'b011011010001010; sin_mem[10'b0101100111] = 15'b010000101111101
    cos_mem[10'b0101101000] = 15'b011011001111101; sin_mem[10'b0101101000] = 15'b010000110010011
    cos_mem[10'b0101101001] = 15'b011011001101111; sin_mem[10'b0101101001] = 15'b010000110101000
    cos_mem[10'b0101101010] = 15'b011011001100010; sin_mem[10'b0101101010] = 15'b010000110111110
    cos_mem[10'b0101101011] = 15'b011011001010101; sin_mem[10'b0101101011] = 15'b010000111010011
    cos_mem[10'b0101101100] = 15'b011011001001000; sin_mem[10'b0101101100] = 15'b010000111101000
    cos_mem[10'b0101101101] = 15'b011011000111010; sin_mem[10'b0101101101] = 15'b010000111111110
    cos_mem[10'b0101101110] = 15'b011011000101101; sin_mem[10'b0101101110] = 15'b010001000010011
    cos_mem[10'b0101101111] = 15'b011011000100000; sin_mem[10'b0101101111] = 15'b010001000101000
    cos_mem[10'b0101110000] = 15'b011011000010010; sin_mem[10'b0101110000] = 15'b010001000111101
    cos_mem[10'b0101110001] = 15'b011011000000101; sin_mem[10'b0101110001] = 15'b010001001010011
    cos_mem[10'b0101110010] = 15'b011010111110111; sin_mem[10'b0101110010] = 15'b010001001101000
    cos_mem[10'b0101110011] = 15'b011010111101010; sin_mem[10'b0101110011] = 15'b010001001111101
    cos_mem[10'b0101110100] = 15'b011010111011100; sin_mem[10'b0101110100] = 15'b010001010010010
    cos_mem[10'b0101110101] = 15'b011010111001110; sin_mem[10'b0101110101] = 15'b010001010100111
    cos_mem[10'b0101110110] = 15'b011010111000001; sin_mem[10'b0101110110] = 15'b010001010111100
    cos_mem[10'b0101110111] = 15'b011010110110011; sin_mem[10'b0101110111] = 15'b010001011010010
    cos_mem[10'b0101111000] = 15'b011010110100101; sin_mem[10'b0101111000] = 15'b010001011100111
    cos_mem[10'b0101111001] = 15'b011010110011000; sin_mem[10'b0101111001] = 15'b010001011111100
    cos_mem[10'b0101111010] = 15'b011010110001010; sin_mem[10'b0101111010] = 15'b010001100010001
    cos_mem[10'b0101111011] = 15'b011010101111100; sin_mem[10'b0101111011] = 15'b010001100100110
    cos_mem[10'b0101111100] = 15'b011010101101110; sin_mem[10'b0101111100] = 15'b010001100111011
    cos_mem[10'b0101111101] = 15'b011010101100001; sin_mem[10'b0101111101] = 15'b010001101010000
    cos_mem[10'b0101111110] = 15'b011010101010011; sin_mem[10'b0101111110] = 15'b010001101100101
    cos_mem[10'b0101111111] = 15'b011010101000101; sin_mem[10'b0101111111] = 15'b010001101111010
    cos_mem[10'b0110000000] = 15'b011010100110111; sin_mem[10'b0110000000] = 15'b010001110001110
    cos_mem[10'b0110000001] = 15'b011010100101001; sin_mem[10'b0110000001] = 15'b010001110100011
    cos_mem[10'b0110000010] = 15'b011010100011011; sin_mem[10'b0110000010] = 15'b010001110111000
    cos_mem[10'b0110000011] = 15'b011010100001101; sin_mem[10'b0110000011] = 15'b010001111001101
    cos_mem[10'b0110000100] = 15'b011010011111111; sin_mem[10'b0110000100] = 15'b010001111100010
    cos_mem[10'b0110000101] = 15'b011010011110001; sin_mem[10'b0110000101] = 15'b010001111110111
    cos_mem[10'b0110000110] = 15'b011010011100010; sin_mem[10'b0110000110] = 15'b010010000001011
    cos_mem[10'b0110000111] = 15'b011010011010100; sin_mem[10'b0110000111] = 15'b010010000100000
    cos_mem[10'b0110001000] = 15'b011010011000110; sin_mem[10'b0110001000] = 15'b010010000110101
    cos_mem[10'b0110001001] = 15'b011010010111000; sin_mem[10'b0110001001] = 15'b010010001001010
    cos_mem[10'b0110001010] = 15'b011010010101010; sin_mem[10'b0110001010] = 15'b010010001011110
    cos_mem[10'b0110001011] = 15'b011010010011011; sin_mem[10'b0110001011] = 15'b010010001110011
    cos_mem[10'b0110001100] = 15'b011010010001101; sin_mem[10'b0110001100] = 15'b010010010001000
    cos_mem[10'b0110001101] = 15'b011010001111111; sin_mem[10'b0110001101] = 15'b010010010011100
    cos_mem[10'b0110001110] = 15'b011010001110000; sin_mem[10'b0110001110] = 15'b010010010110001
    cos_mem[10'b0110001111] = 15'b011010001100010; sin_mem[10'b0110001111] = 15'b010010011000101
    cos_mem[10'b0110010000] = 15'b011010001010011; sin_mem[10'b0110010000] = 15'b010010011011010
    cos_mem[10'b0110010001] = 15'b011010001000101; sin_mem[10'b0110010001] = 15'b010010011101111
    cos_mem[10'b0110010010] = 15'b011010000110110; sin_mem[10'b0110010010] = 15'b010010100000011
    cos_mem[10'b0110010011] = 15'b011010000101000; sin_mem[10'b0110010011] = 15'b010010100011000
    cos_mem[10'b0110010100] = 15'b011010000011001; sin_mem[10'b0110010100] = 15'b010010100101100
    cos_mem[10'b0110010101] = 15'b011010000001011; sin_mem[10'b0110010101] = 15'b010010101000001
    cos_mem[10'b0110010110] = 15'b011001111111100; sin_mem[10'b0110010110] = 15'b010010101010101
    cos_mem[10'b0110010111] = 15'b011001111101101; sin_mem[10'b0110010111] = 15'b010010101101001
    cos_mem[10'b0110011000] = 15'b011001111011111; sin_mem[10'b0110011000] = 15'b010010101111110
    cos_mem[10'b0110011001] = 15'b011001111010000; sin_mem[10'b0110011001] = 15'b010010110010010
    cos_mem[10'b0110011010] = 15'b011001111000001; sin_mem[10'b0110011010] = 15'b010010110100110
    cos_mem[10'b0110011011] = 15'b011001110110010; sin_mem[10'b0110011011] = 15'b010010110111011
    cos_mem[10'b0110011100] = 15'b011001110100011; sin_mem[10'b0110011100] = 15'b010010111001111
    cos_mem[10'b0110011101] = 15'b011001110010101; sin_mem[10'b0110011101] = 15'b010010111100011
    cos_mem[10'b0110011110] = 15'b011001110000110; sin_mem[10'b0110011110] = 15'b010010111111000
    cos_mem[10'b0110011111] = 15'b011001101110111; sin_mem[10'b0110011111] = 15'b010011000001100
    cos_mem[10'b0110100000] = 15'b011001101101000; sin_mem[10'b0110100000] = 15'b010011000100000
    cos_mem[10'b0110100001] = 15'b011001101011001; sin_mem[10'b0110100001] = 15'b010011000110100
    cos_mem[10'b0110100010] = 15'b011001101001010; sin_mem[10'b0110100010] = 15'b010011001001000
    cos_mem[10'b0110100011] = 15'b011001100111011; sin_mem[10'b0110100011] = 15'b010011001011100
    cos_mem[10'b0110100100] = 15'b011001100101100; sin_mem[10'b0110100100] = 15'b010011001110001
    cos_mem[10'b0110100101] = 15'b011001100011101; sin_mem[10'b0110100101] = 15'b010011010000101
    cos_mem[10'b0110100110] = 15'b011001100001101; sin_mem[10'b0110100110] = 15'b010011010011001
    cos_mem[10'b0110100111] = 15'b011001011111110; sin_mem[10'b0110100111] = 15'b010011010101101
    cos_mem[10'b0110101000] = 15'b011001011101111; sin_mem[10'b0110101000] = 15'b010011011000001
    cos_mem[10'b0110101001] = 15'b011001011100000; sin_mem[10'b0110101001] = 15'b010011011010101
    cos_mem[10'b0110101010] = 15'b011001011010000; sin_mem[10'b0110101010] = 15'b010011011101001
    cos_mem[10'b0110101011] = 15'b011001011000001; sin_mem[10'b0110101011] = 15'b010011011111101
    cos_mem[10'b0110101100] = 15'b011001010110010; sin_mem[10'b0110101100] = 15'b010011100010001
    cos_mem[10'b0110101101] = 15'b011001010100011; sin_mem[10'b0110101101] = 15'b010011100100100
    cos_mem[10'b0110101110] = 15'b011001010010011; sin_mem[10'b0110101110] = 15'b010011100111000
    cos_mem[10'b0110101111] = 15'b011001010000100; sin_mem[10'b0110101111] = 15'b010011101001100
    cos_mem[10'b0110110000] = 15'b011001001110100; sin_mem[10'b0110110000] = 15'b010011101100000
    cos_mem[10'b0110110001] = 15'b011001001100101; sin_mem[10'b0110110001] = 15'b010011101110100
    cos_mem[10'b0110110010] = 15'b011001001010101; sin_mem[10'b0110110010] = 15'b010011110001000
    cos_mem[10'b0110110011] = 15'b011001001000110; sin_mem[10'b0110110011] = 15'b010011110011011
    cos_mem[10'b0110110100] = 15'b011001000110110; sin_mem[10'b0110110100] = 15'b010011110101111
    cos_mem[10'b0110110101] = 15'b011001000100111; sin_mem[10'b0110110101] = 15'b010011111000011
    cos_mem[10'b0110110110] = 15'b011001000010111; sin_mem[10'b0110110110] = 15'b010011111010110
    cos_mem[10'b0110110111] = 15'b011001000000111; sin_mem[10'b0110110111] = 15'b010011111101010
    cos_mem[10'b0110111000] = 15'b011000111111000; sin_mem[10'b0110111000] = 15'b010011111111110
    cos_mem[10'b0110111001] = 15'b011000111101000; sin_mem[10'b0110111001] = 15'b010100000010001
    cos_mem[10'b0110111010] = 15'b011000111011000; sin_mem[10'b0110111010] = 15'b010100000100101
    cos_mem[10'b0110111011] = 15'b011000111001000; sin_mem[10'b0110111011] = 15'b010100000111000
    cos_mem[10'b0110111100] = 15'b011000110111001; sin_mem[10'b0110111100] = 15'b010100001001100
    cos_mem[10'b0110111101] = 15'b011000110101001; sin_mem[10'b0110111101] = 15'b010100001100000
    cos_mem[10'b0110111110] = 15'b011000110011001; sin_mem[10'b0110111110] = 15'b010100001110011
    cos_mem[10'b0110111111] = 15'b011000110001001; sin_mem[10'b0110111111] = 15'b010100010000110
    cos_mem[10'b0111000000] = 15'b011000101111001; sin_mem[10'b0111000000] = 15'b010100010011010
    cos_mem[10'b0111000001] = 15'b011000101101001; sin_mem[10'b0111000001] = 15'b010100010101101
    cos_mem[10'b0111000010] = 15'b011000101011001; sin_mem[10'b0111000010] = 15'b010100011000001
    cos_mem[10'b0111000011] = 15'b011000101001001; sin_mem[10'b0111000011] = 15'b010100011010100
    cos_mem[10'b0111000100] = 15'b011000100111001; sin_mem[10'b0111000100] = 15'b010100011100111
    cos_mem[10'b0111000101] = 15'b011000100101001; sin_mem[10'b0111000101] = 15'b010100011111011
    cos_mem[10'b0111000110] = 15'b011000100011001; sin_mem[10'b0111000110] = 15'b010100100001110
    cos_mem[10'b0111000111] = 15'b011000100001001; sin_mem[10'b0111000111] = 15'b010100100100001
    cos_mem[10'b0111001000] = 15'b011000011111001; sin_mem[10'b0111001000] = 15'b010100100110101
    cos_mem[10'b0111001001] = 15'b011000011101000; sin_mem[10'b0111001001] = 15'b010100101001000
    cos_mem[10'b0111001010] = 15'b011000011011000; sin_mem[10'b0111001010] = 15'b010100101011011
    cos_mem[10'b0111001011] = 15'b011000011001000; sin_mem[10'b0111001011] = 15'b010100101101110
    cos_mem[10'b0111001100] = 15'b011000010111000; sin_mem[10'b0111001100] = 15'b010100110000001
    cos_mem[10'b0111001101] = 15'b011000010100111; sin_mem[10'b0111001101] = 15'b010100110010100
    cos_mem[10'b0111001110] = 15'b011000010010111; sin_mem[10'b0111001110] = 15'b010100110100111
    cos_mem[10'b0111001111] = 15'b011000010000111; sin_mem[10'b0111001111] = 15'b010100110111011
    cos_mem[10'b0111010000] = 15'b011000001110110; sin_mem[10'b0111010000] = 15'b010100111001110
    cos_mem[10'b0111010001] = 15'b011000001100110; sin_mem[10'b0111010001] = 15'b010100111100001
    cos_mem[10'b0111010010] = 15'b011000001010101; sin_mem[10'b0111010010] = 15'b010100111110100
    cos_mem[10'b0111010011] = 15'b011000001000101; sin_mem[10'b0111010011] = 15'b010101000000111
    cos_mem[10'b0111010100] = 15'b011000000110100; sin_mem[10'b0111010100] = 15'b010101000011010
    cos_mem[10'b0111010101] = 15'b011000000100100; sin_mem[10'b0111010101] = 15'b010101000101100
    cos_mem[10'b0111010110] = 15'b011000000010011; sin_mem[10'b0111010110] = 15'b010101000111111
    cos_mem[10'b0111010111] = 15'b011000000000010; sin_mem[10'b0111010111] = 15'b010101001010010
    cos_mem[10'b0111011000] = 15'b010111111110010; sin_mem[10'b0111011000] = 15'b010101001100101
    cos_mem[10'b0111011001] = 15'b010111111100001; sin_mem[10'b0111011001] = 15'b010101001111000
    cos_mem[10'b0111011010] = 15'b010111111010000; sin_mem[10'b0111011010] = 15'b010101010001011
    cos_mem[10'b0111011011] = 15'b010111111000000; sin_mem[10'b0111011011] = 15'b010101010011101
    cos_mem[10'b0111011100] = 15'b010111110101111; sin_mem[10'b0111011100] = 15'b010101010110000
    cos_mem[10'b0111011101] = 15'b010111110011110; sin_mem[10'b0111011101] = 15'b010101011000011
    cos_mem[10'b0111011110] = 15'b010111110001101; sin_mem[10'b0111011110] = 15'b010101011010110
    cos_mem[10'b0111011111] = 15'b010111101111101; sin_mem[10'b0111011111] = 15'b010101011101000
    cos_mem[10'b0111100000] = 15'b010111101101100; sin_mem[10'b0111100000] = 15'b010101011111011
    cos_mem[10'b0111100001] = 15'b010111101011011; sin_mem[10'b0111100001] = 15'b010101100001101
    cos_mem[10'b0111100010] = 15'b010111101001010; sin_mem[10'b0111100010] = 15'b010101100100000
    cos_mem[10'b0111100011] = 15'b010111100111001; sin_mem[10'b0111100011] = 15'b010101100110011
    cos_mem[10'b0111100100] = 15'b010111100101000; sin_mem[10'b0111100100] = 15'b010101101000101
    cos_mem[10'b0111100101] = 15'b010111100010111; sin_mem[10'b0111100101] = 15'b010101101011000
    cos_mem[10'b0111100110] = 15'b010111100000110; sin_mem[10'b0111100110] = 15'b010101101101010
    cos_mem[10'b0111100111] = 15'b010111011110101; sin_mem[10'b0111100111] = 15'b010101101111101
    cos_mem[10'b0111101000] = 15'b010111011100100; sin_mem[10'b0111101000] = 15'b010101110001111
    cos_mem[10'b0111101001] = 15'b010111011010011; sin_mem[10'b0111101001] = 15'b010101110100001
    cos_mem[10'b0111101010] = 15'b010111011000010; sin_mem[10'b0111101010] = 15'b010101110110100
    cos_mem[10'b0111101011] = 15'b010111010110000; sin_mem[10'b0111101011] = 15'b010101111000110
    cos_mem[10'b0111101100] = 15'b010111010011111; sin_mem[10'b0111101100] = 15'b010101111011000
    cos_mem[10'b0111101101] = 15'b010111010001110; sin_mem[10'b0111101101] = 15'b010101111101011
    cos_mem[10'b0111101110] = 15'b010111001111101; sin_mem[10'b0111101110] = 15'b010101111111101
    cos_mem[10'b0111101111] = 15'b010111001101011; sin_mem[10'b0111101111] = 15'b010110000001111
    cos_mem[10'b0111110000] = 15'b010111001011010; sin_mem[10'b0111110000] = 15'b010110000100001
    cos_mem[10'b0111110001] = 15'b010111001001001; sin_mem[10'b0111110001] = 15'b010110000110100
//cut here----------------------------------------------------------------------------------------------    
    cos_mem[10'b0111110010] = 15'b010111000110111; sin_mem[10'b0111110010] = 15'b010110001000110
    cos_mem[10'b0111110011] = 15'b010111000100110; sin_mem[10'b0111110011] = 15'b010110001011000
    cos_mem[10'b0111110100] = 15'b010111000010101; sin_mem[10'b0111110100] = 15'b010110001101010
    cos_mem[10'b0111110101] = 15'b010111000000011; sin_mem[10'b0111110101] = 15'b010110001111100
    cos_mem[10'b0111110110] = 15'b010110111110010; sin_mem[10'b0111110110] = 15'b010110010001110
    cos_mem[10'b0111110111] = 15'b010110111100000; sin_mem[10'b0111110111] = 15'b010110010100000
    cos_mem[10'b0111111000] = 15'b010110111001111; sin_mem[10'b0111111000] = 15'b010110010110010
    cos_mem[10'b0111111001] = 15'b010110110111101; sin_mem[10'b0111111001] = 15'b010110011000100
    cos_mem[10'b0111111010] = 15'b010110110101011; sin_mem[10'b0111111010] = 15'b010110011010110
    cos_mem[10'b0111111011] = 15'b010110110011010; sin_mem[10'b0111111011] = 15'b010110011101000
    cos_mem[10'b0111111100] = 15'b010110110001000; sin_mem[10'b0111111100] = 15'b010110011111010
    cos_mem[10'b0111111101] = 15'b010110101110110; sin_mem[10'b0111111101] = 15'b010110100001100
    cos_mem[10'b0111111110] = 15'b010110101100101; sin_mem[10'b0111111110] = 15'b010110100011110
    cos_mem[10'b0111111111] = 15'b010110101010011; sin_mem[10'b0111111111] = 15'b010110100101111
    cos_mem[10'b1000000000] = 15'b010110101000001; sin_mem[10'b1000000000] = 15'b010110101000001
end

always @(angle or cos_en) begin
    //cos/sin selection for output
    if (cos_en == 1'b1)
        //compute cos(angle)
        angle_output = angle;
    else
        //compute sin(angle) = cos (pi/2 - angle)
        angle_output = 11'b100_0000_0000 - angle;

    //choose cos/sin mem bank
    case (angle_output[11:9])
        3'b000: begin //0 - 45
            angle_mem_full = angle_output;
            select_cos_mem = 1'b1;
            select_positive = 1'b1;
        end
        3'b001: begin //45 - 90
            angle_mem_full = 12'h400 - angle_output;
            select_cos_mem = 1'b0;
            select_positive = 1'b1;
        end
        3'b010: begin //90 - 135
            angle_mem_full = angle_output[9:0] - 12'h400;
            select_cos_mem = 1'b0;
            select_positive = 1'b0;
        end
        3'b011: begin //135 - 180
            angle_mem_full = 12'h800 - angle_output;
            select_cos_mem = 1'b1;
            select_positive = 1'b0;
        end
        3'b100: begin //180 - 225
            angle_mem_full = angle_output - 12'h800;
            select_cos_mem = 1'b1;
            select_positive = 1'b0;
        end
        3'b101: begin //225 - 270
            angle_mem_full = 12'hC00 - angle_output;
            select_cos_mem = 1'b0;
            select_positive = 1'b0;
        end
        3'b110: begin //270 - 315
            angle_mem_full = angle_output - 12'hC00;
            select_cos_mem = 1'b0;
            select_positive = 1'b1;
        end
        3'b111: begin //315 - 360
            angle_mem_full = 13'h1000 - angle_output;
            select_cos_mem = 1'b1;
            select_positive = 1'b1;
        end
    endcase

    //read memory
    angle_mem = angle_output[10:0];
    if (select_cos_mem == 1'b1) begin
        if (select_positive) begin
            mem_val = cos_mem[angle_mem];
        end else begin
            mem_val = -cos_mem[angle_mem];
        end
    end else begin
        if (select_positive) begin
            mem_val = sin_mem[angle_mem];
        end else begin
            mem_val = -sin_mem[angle_mem];
        end
    end

    //exception (when need to return +1.0)
    except = (angle_mem == 10'b00_0000_0000);
    except = except || (angle_mem == 10'b00_0000_0001);
    except = except || (angle_mem == 10'b00_0000_0010);
    except = except || (angle_mem == 10'b00_0000_0011);
    except = except || (angle_mem == 10'b00_0000_0100);
    except = except || (angle_mem == 10'b00_0000_0101);
    //except only work for cos bank near angle 0
    except = except & select_cos_mem;

    //make output
    result = {mem_val[14], mem_val[14] | except, mem_val[13:0]};
end

endmodule