//fixed to float

`timescale 1ns/10ps

module fxfl(
  input [6:0] fx,
  output reg [3:0] m,
  output reg [3:0] e
);

always @(fx)
  casez (fx)
    7'b0000000: {m,e} = 8'b00000000;
  //positive numbers
    7'b0000001: {m,e} = 8'b01001011;        //0100 * 2^(-5)
    7'b000001?: {m,e} = {fx[2:0],5'b01100}; //01x0 * 2^(-4)
    7'b00001??: {m,e} = {fx[3:0],4'b1101};  //01xx * 2^(-3)
    7'b0001???: {m,e} = {fx[4:1],4'b1110};  //01xx * 2^(-2)
    7'b001????: {m,e} = {fx[5:2],4'b1111};  //01xx * 2^(-1)
    7'b01?????: {m,e} = {fx[6:3],4'b0000};  //01xx * 2^( 0)
  //negative numbers
    7'b1111111: {m,e} = 8'b10001010;        //1000 * 2^(-6)
    7'b1111110: {m,e} = 8'b10001011;        //1000 * 2^(-5)
    7'b11111??: {m,e} = {fx[2:0],5'b01100}; //1xx0 * 2^(-4)
    7'b1111???: {m,e} = {fx[3:0],4'b1101};  //1xxx * 2^(-3)
    7'b111????: {m,e} = {fx[4:1],4'b1110};  //1xxx * 2^(-2)
    7'b11?????: {m,e} = {fx[5:2],4'b1111};  //1xxx * 2^(-1)
    7'b1??????: {m,e} = {fx[6:3],4'b0000};  //1xxx * 2^( 0)
    default: {m,e} = 8'h0f;
  endcase

endmodule
