//HW2 P2
//

`timescale 1ns/10ps

module mult8x8 (
    input reg [7:0] a,
    input reg [7:0] b,
    output reg [15:0] out
);

//stage 1. encoding
    reg [7:0] pp0,pp1,pp2,pp3,pp4,pp5,pp6,pp7;
    always @(a or b) begin
        pp0 = {~a[7],a[6:0]} & {b[0], b[0], b[0], b[0], b[0], b[0], b[0], b[0]};
        pp1 = {~a[7],a[6:0]} & {b[1], b[1], b[1], b[1], b[1], b[1], b[1], b[1]};
        pp2 = {~a[7],a[6:0]} & {b[2], b[2], b[2], b[2], b[2], b[2], b[2], b[2]};
        pp3 = {~a[7],a[6:0]} & {b[3], b[3], b[3], b[3], b[3], b[3], b[3], b[3]};
        pp4 = {~a[7],a[6:0]} & {b[4], b[4], b[4], b[4], b[4], b[4], b[4], b[4]};
        pp5 = {~a[7],a[6:0]} & {b[5], b[5], b[5], b[5], b[5], b[5], b[5], b[5]};
        pp6 = {~a[7],a[6:0]} & {b[6], b[6], b[6], b[6], b[6], b[6], b[6], b[6]};
        pp7 = {~a[7],a[6:0]} & {b[7], b[7], b[7], b[7], b[7], b[7], b[7], b[7]};
    end

//stage 2. CSA
/*  0         -.......
    1        -.......
    2       -.......
    3      -.......
    4     -.......
    5    -.......
    6   -.......
    7  -.......
    8 111111111
    9 11111111
    a 1111111
    b 111111
    c 11111
    d 1111
    e 111
    f 11
      ================
    0         -.......
    1        -.......
    2       -.......
    3      -.......
    4     -.......
    5    -.......
    6   -.......
    7  -.......
    8 100000001
      ================
*/

      
endmodule
